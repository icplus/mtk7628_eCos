# ====================================================================
#
#      openssl.cdl
#
#      openssl configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      andrew Lunn
# Original data:  andrew Lunn
# Contributors:   Andrew Lunn
# Date:           2001-05-22
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_OPENSSL {
    display       "OpenSSL"
    parent        CYGPKG_NET
#    doc           doc/index.html
    include_dir   openssl
    requires      CYGPKG_IO
    requires      CYGPKG_LIBC
    requires      CYGPKG_ERROR
    requires      CYGPKG_NET
# RAND requires that there is at least one message digest algorithm
    requires      { (CYGPKG_OPENSSL_SHA && CYGPKG_OPENSSL_SHA1) || 
                    CYGPKG_OPENSSL_MD5 || 
                    (CYGPKG_OPENSSL_MDC2 && CYGPKG_OPENSSL_DES) ||
                    (CYGPKG_OPENSSL_MD2) }
# x_name appears to be broken without buffer
    requires      CYGPKG_OPENSSL_BUFFER  
# txt_db appears to be broken without BIO
    requires      CYGPKG_OPENSSL_BIO
    description   "Port of the OpenSSL library."

    compile					\
        crypto/asn1/a_object.c  \
        crypto/asn1/a_bitstr.c  \
        crypto/asn1/a_utctm.c   \
        crypto/asn1/a_gentm.c   \
        crypto/asn1/a_time.c    \
        crypto/asn1/a_int.c     \
        crypto/asn1/a_octet.c   \
        crypto/asn1/a_null.c    \
        crypto/asn1/a_print.c   \
        crypto/asn1/a_type.c    \
        crypto/asn1/a_set.c     \
        crypto/asn1/a_dup.c     \
        crypto/asn1/a_d2i_fp.c  \
        crypto/asn1/a_i2d_fp.c  \
        crypto/asn1/a_bmp.c     \
        crypto/asn1/a_enum.c    \
        crypto/asn1/a_vis.c     \
        crypto/asn1/a_utf8.c    \
        crypto/asn1/a_sign.c    \
        crypto/asn1/a_digest.c  \
        crypto/asn1/a_verify.c  \
        crypto/asn1/a_mbstr.c   \
        crypto/asn1/a_strex.c   \
        crypto/asn1/x_algor.c   \
        crypto/asn1/x_val.c     \
        crypto/asn1/x_pubkey.c  \
        crypto/asn1/x_sig.c     \
        crypto/asn1/x_req.c     \
        crypto/asn1/x_attrib.c  \
        crypto/asn1/x_name.c    \
        crypto/asn1/x_cinf.c    \
        crypto/asn1/x_x509.c    \
        crypto/asn1/x_x509a.c   \
        crypto/asn1/x_crl.c     \
        crypto/asn1/x_info.c    \
        crypto/asn1/x_spki.c    \
        crypto/asn1/nsseq.c     \
        crypto/asn1/d2i_r_pr.c  \
        crypto/asn1/i2d_r_pr.c  \
        crypto/asn1/d2i_r_pu.c  \
        crypto/asn1/i2d_r_pu.c  \
        crypto/asn1/d2i_s_pr.c  \
        crypto/asn1/i2d_s_pr.c  \
        crypto/asn1/d2i_s_pu.c  \
        crypto/asn1/i2d_s_pu.c  \
        crypto/asn1/d2i_pu.c    \
        crypto/asn1/d2i_pr.c    \
        crypto/asn1/i2d_pu.c    \
        crypto/asn1/i2d_pr.c    \
        crypto/asn1/t_req.c     \
        crypto/asn1/t_x509.c    \
        crypto/asn1/t_x509a.c   \
        crypto/asn1/t_crl.c     \
        crypto/asn1/t_pkey.c    \
        crypto/asn1/t_spki.c    \
        crypto/asn1/t_bitst.c   \
        crypto/asn1/p7_i_s.c    \
        crypto/asn1/p7_signi.c  \
        crypto/asn1/p7_signd.c  \
        crypto/asn1/p7_recip.c  \
        crypto/asn1/p7_enc_c.c  \
        crypto/asn1/p7_evp.c    \
        crypto/asn1/p7_dgst.c   \
        crypto/asn1/p7_s_e.c    \
        crypto/asn1/p7_enc.c    \
        crypto/asn1/p7_lib.c    \
        crypto/asn1/f_int.c     \
        crypto/asn1/f_string.c  \
        crypto/asn1/i2d_dhp.c   \
        crypto/asn1/i2d_dsap.c  \
        crypto/asn1/d2i_dhp.c   \
        crypto/asn1/d2i_dsap.c  \
        crypto/asn1/n_pkey.c    \
        crypto/asn1/f_enum.c    \
        crypto/asn1/a_hdr.c     \
        crypto/asn1/x_pkey.c    \
        crypto/asn1/a_bool.c    \
        crypto/asn1/x_exten.c   \
        crypto/asn1/asn1_par.c  \
        crypto/asn1/asn1_lib.c  \
        crypto/asn1/asn1_err.c  \
        crypto/asn1/a_meth.c    \
        crypto/asn1/a_bytes.c   \
        crypto/asn1/a_strnid.c  \
        crypto/asn1/evp_asn1.c  \
        crypto/asn1/asn_pack.c  \
        crypto/asn1/p5_pbe.c    \
        crypto/asn1/p5_pbev2.c  \
        crypto/asn1/p8_pkey.c   \
        crypto/bn/bn_add.c      \
        crypto/bn/bn_div.c      \
        crypto/bn/bn_exp.c      \
        crypto/bn/bn_lib.c      \
        crypto/bn/bn_ctx.c      \
        crypto/bn/bn_mul.c      \
        crypto/bn/bn_print.c    \
        crypto/bn/bn_rand.c     \
        crypto/bn/bn_shift.c    \
        crypto/bn/bn_word.c     \
        crypto/bn/bn_blind.c    \
        crypto/bn/bn_gcd.c      \
        crypto/bn/bn_prime.c    \
        crypto/bn/bn_err.c      \
        crypto/bn/bn_sqr.c      \
        crypto/bn/bn_asm.c      \
        crypto/bn/bn_recp.c     \
        crypto/bn/bn_mont.c     \
        crypto/bn/bn_mpi.c      \
        crypto/bn/bn_exp2.c     \
        crypto/evp/encode.c     \
        crypto/evp/digest.c     \
        crypto/evp/evp_enc.c    \
        crypto/evp/evp_key.c    \
        crypto/evp/e_des.c      \
        crypto/evp/e_bf.c       \
        crypto/evp/e_idea.c     \
        crypto/evp/e_des3.c     \
        crypto/evp/e_rc4.c      \
        crypto/evp/names.c      \
        crypto/evp/e_xcbc_d.c   \
        crypto/evp/e_rc2.c      \
        crypto/evp/e_cast.c     \
        crypto/evp/e_rc5.c      \
        crypto/evp/m_null.c     \
        crypto/evp/m_md2.c      \
        crypto/evp/m_md4.c      \
        crypto/evp/m_md5.c      \
        crypto/evp/m_sha.c      \
        crypto/evp/m_sha1.c     \
        crypto/evp/m_dss.c      \
        crypto/evp/m_dss1.c     \
        crypto/evp/m_mdc2.c     \
        crypto/evp/m_ripemd.c   \
        crypto/evp/p_open.c     \
        crypto/evp/p_seal.c     \
        crypto/evp/p_sign.c     \
        crypto/evp/p_verify.c   \
        crypto/evp/p_lib.c      \
        crypto/evp/p_enc.c      \
        crypto/evp/p_dec.c      \
        crypto/evp/bio_md.c     \
        crypto/evp/bio_b64.c    \
        crypto/evp/bio_enc.c    \
        crypto/evp/evp_err.c    \
        crypto/evp/e_null.c     \
        crypto/evp/c_all.c      \
        crypto/evp/c_allc.c     \
        crypto/evp/c_alld.c     \
        crypto/evp/evp_lib.c    \
        crypto/evp/bio_ok.c     \
        crypto/evp/evp_pkey.c   \
        crypto/evp/evp_pbe.c    \
        crypto/evp/p5_crpt.c    \
        crypto/evp/p5_crpt2.c   \
        crypto/hmac/hmac.c      \
        crypto/lhash/lhash.c    \
        crypto/lhash/lh_stats.c \
        crypto/objects/o_names.c \
        crypto/objects/obj_dat.c \
        crypto/objects/obj_lib.c \
        crypto/objects/obj_err.c \
        crypto/pem/pem_sign.c    \
        crypto/pem/pem_seal.c   \
        crypto/pem/pem_info.c   \
        crypto/pem/pem_lib.c    \
        crypto/pem/pem_all.c    \
        crypto/pem/pem_err.c    \
        crypto/pkcs7/pk7_lib.c  \
        crypto/pkcs7/pkcs7err.c \
        crypto/pkcs7/pk7_doit.c \
        crypto/pkcs7/pk7_smime.c \
        crypto/pkcs7/pk7_attr.c  \
        crypto/pkcs7/pk7_mime.c  \
        crypto/pkcs12/p12_add.c  \
        crypto/pkcs12/p12_attr.c \
        crypto/pkcs12/p12_bags.c \
        crypto/pkcs12/p12_crpt.c \
        crypto/pkcs12/p12_crt.c  \
        crypto/pkcs12/p12_decr.c \
        crypto/pkcs12/p12_init.c \
        crypto/pkcs12/p12_key.c  \
        crypto/pkcs12/p12_kiss.c \
        crypto/pkcs12/p12_lib.c  \
        crypto/pkcs12/p12_mac.c  \
        crypto/pkcs12/p12_mutl.c \
        crypto/pkcs12/p12_sbag.c \
        crypto/pkcs12/p12_utl.c  \
        crypto/pkcs12/p12_npas.c \
        crypto/pkcs12/pk12err.c \
        crypto/rand/md_rand.c   \
        crypto/rand/randfile.c  \
        crypto/rand/rand_lib.c  \
        crypto/rand/rand_err.c  \
        crypto/rand/rand_egd.c  \
        crypto/rand/rand_win.c  \
        crypto/stack/stack.c    \
        crypto/txt_db/txt_db.c  \
        crypto/x509/x509_def.c  \
        crypto/x509/x509_d2.c   \
        crypto/x509/x509_r2x.c  \
        crypto/x509/x509_cmp.c  \
        crypto/x509/x509_obj.c  \
        crypto/x509/x509_req.c  \
        crypto/x509/x509spki.c  \
        crypto/x509/x509_vfy.c  \
        crypto/x509/x509_set.c  \
        crypto/x509/x509rset.c  \
        crypto/x509/x509_err.c  \
        crypto/x509/x509name.c  \
        crypto/x509/x509_v3.c   \
        crypto/x509/x509_ext.c  \
        crypto/x509/x509_att.c  \
        crypto/x509/x509type.c  \
        crypto/x509/x509_lu.c   \
        crypto/x509/x_all.c     \
        crypto/x509/x509_txt.c  \
        crypto/x509/x509_trs.c  \
        crypto/x509/by_file.c   \
        crypto/x509/by_dir.c    \
        crypto/x509v3/v3_bcons.c \
        crypto/x509v3/v3_bitst.c \
        crypto/x509v3/v3_conf.c  \
        crypto/x509v3/v3_extku.c \
        crypto/x509v3/v3_ia5.c  \
        crypto/x509v3/v3_lib.c  \
        crypto/x509v3/v3_prn.c  \
        crypto/x509v3/v3_utl.c  \
        crypto/x509v3/v3err.c   \
        crypto/x509v3/v3_genn.c \
        crypto/x509v3/v3_alt.c  \
        crypto/x509v3/v3_skey.c \
        crypto/x509v3/v3_akey.c \
        crypto/x509v3/v3_pku.c  \
        crypto/x509v3/v3_int.c  \
        crypto/x509v3/v3_enum.c \
        crypto/x509v3/v3_sxnet.c \
        crypto/x509v3/v3_cpols.c \
        crypto/x509v3/v3_crld.c  \
        crypto/x509v3/v3_purp.c \
        crypto/x509v3/v3_info.c \
        crypto/conf/conf_err.c  \
        crypto/conf/conf_lib.c  \
        crypto/conf/conf_api.c  \
        crypto/conf/conf_def.c  \
        crypto/err/err_all.c    \
        crypto/err/err_prn.c    \
        crypto/err/err.c        \
        crypto/cryptlib.c       \
        crypto/mem.c            \
        crypto/mem_dbg.c        \
        crypto/cversion.c       \
        crypto/ex_data.c        \
        crypto/cpt_err.c        \
        crypto/ebcdic.c         \
        crypto/uid.c            

    cdl_component CYGPKG_OPENSSL_IDEA {
        display       "IDEA encryption algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 0
        description   "
             Implements the IDEA encryption Algorith. Disabled by default

             NOTE: 

             The IDEA algorithm is patented by Ascom in Austria, France, 
             Germany, Italy, Japan, Netherlands, Spain, Sweden, Switzerland, 
             UK and the USA.  They should be contacted if that algorithm is 
             to be used, their web page is http://www.ascom.ch."

        compile        crypto/idea/i_cbc.c     \
                       crypto/idea/i_cfb64.c   \
                       crypto/idea/i_ofb64.c   \
                       crypto/idea/i_ecb.c     \
                       crypto/idea/i_skey.c    
    }
    cdl_option CYGPKG_OPENSSL_IDEA_TESTS {
        display "OpenSSL IDEA tests"
        flavor  data
        no_define
        calculated { " tests/ideatest.c" }
        description   "
            This option specifies the test for the idea algorithm"
    }
    cdl_component CYGPKG_OPENSSL_RC5 {
        display       "RC5 encryption algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 0
        description   "
             Implements the RC5 encryption Algorith. Disabled by default

             NOTE: 

             RSA Data Security holds software patents on the RSA and
             RC5 algorithms.  If their ciphers are used used inside
             the USA (and Japan?), you must contact RSA Data Security
             for licencing conditions.  Their web page is http://www.rsa.com"

        compile       crypto/rc5/rc5_skey.c   \
                      crypto/rc5/rc5_ecb.c    \
                      crypto/rc5/rc5_enc.c    \
                      crypto/rc5/rc5cfb64.c   \
                      crypto/rc5/rc5ofb64.c   
     }
     cdl_option CYGPKG_OPENSSL_RC5_TESTS {
         display "OpenSSL RC5 tests"
         flavor  data
         no_define
         calculated { 
            " tests/rc5test.c"
         }
         description   "
             This option specifies the test for the RC5 algorithm"
    }
    cdl_component CYGPKG_OPENSSL_RSA {
        display       "RSA encryption algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 0
        description   "
             Implements the RSA encryption Algorith. Disabled by default

             NOTE: 

             RSA Data Security holds software patents on the RSA and
             RC5 algorithms.  If their ciphers are used used inside
             the USA (and Japan?), you must contact RSA Data Security
             for licencing conditions.  Their web page is http://www.rsa.com"

        compile        crypto/rsa/rsa_eay.c    \
                       crypto/rsa/rsa_gen.c    \
                       crypto/rsa/rsa_lib.c    \
                       crypto/rsa/rsa_sign.c   \
                       crypto/rsa/rsa_saos.c   \
                       crypto/rsa/rsa_err.c    \
                       crypto/rsa/rsa_pk1.c    \
                       crypto/rsa/rsa_ssl.c    \
                       crypto/rsa/rsa_none.c   \
                       crypto/rsa/rsa_oaep.c   \
                       crypto/rsa/rsa_null.c
    }    
    cdl_option CYGPKG_OPENSSL_RSA_TESTS {
         display "OpenSSL RSA tests"
         flavor  data
         no_define
         default_value { " tests/rsa_test.c"}
         description   "
                 This option specifies the test for the RSA algorithm"
    }
    cdl_component CYGPKG_OPENSSL_MD2 {
        display       "MD2 algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the MD2 Algorithm."

        compile        crypto/md2/md2_dgst.c   \
                       crypto/md2/md2_one.c   
    }                
    cdl_option CYGPKG_OPENSSL_MD2_TESTS {
        display "OpenSSL MD2 tests"
        flavor  data
        no_define
        calculated { 
           " tests/md2test.c"
        }
        description   "
            This option specifies the test for the md2 algorithm"
    }
    cdl_component CYGPKG_OPENSSL_MD4 {
        display       "MD4 algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the MD4 Algorith."

        compile        crypto/md4/md4_dgst.c   \
                       crypto/md4/md4_one.c   
    }                  
    cdl_option CYGPKG_OPENSSL_MD4_TESTS {
        display "OpenSSL MD4 tests"
        flavor  data
        no_define
        calculated { 
           " tests/md4test.c"
        }
        description   "
            This option specifies the test for the md4 algorithm"
    }
    cdl_component CYGPKG_OPENSSL_MD5 {
        display       "MD5 algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the MD5 Algorith."

        compile        crypto/md5/md5_dgst.c   \
                       crypto/md5/md5_one.c   
    }                
    cdl_option CYGPKG_OPENSSL_MD5_TESTS {
        display "OpenSSL MD5 tests"
        flavor  data
        no_define
        calculated { 
           " tests/md5test.c"
        }
        description   "
             This option specifies the test for the md5 algorithm"
    }
    cdl_component CYGPKG_OPENSSL_SHA {
        display       "SHA algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the SHA Algorith."

        compile        crypto/sha/sha_dgst.c   \
                       crypto/sha/sha_one.c   
    }                
    cdl_option CYGPKG_OPENSSL_SHA_TESTS {
        display "OpenSSL SHA tests"
        flavor  data
        no_define
        calculated { 
           " tests/shatest.c"
        }
        description   "
            This option specifies the test for the sha algorithm"
    }
    cdl_component CYGPKG_OPENSSL_SHA1 {
        display       "SHA1 algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        requires      CYGPKG_OPENSSL_SHA
        default_value 1
        description   "
             Implements the SHA1 Algorith."

        compile        crypto/sha/sha1dgst.c   \
                       crypto/sha/sha1_one.c   
    }                
    cdl_option CYGPKG_OPENSSL_SHA1_TESTS {
        display "OpenSSL SHA1 tests"
        flavor  data
        no_define
        calculated { 
           " tests/sha1test.c"
        }
        description   "
            This option specifies the test for the sha1 algorithm"
    }
    cdl_component CYGPKG_OPENSSL_RMD160 {
        display       "RMD 160 algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the RMD 160 Algorith."

        compile        crypto/ripemd/rmd_dgst.c   \
                       crypto/ripemd/rmd_one.c   
    }            
    cdl_option CYGPKG_OPENSSL_RMD160_TESTS {
        display "OpenSSL RMD160 tests"
        flavor  data
        no_define
        calculated { 
           " tests/rmdtest.c"
        }
        description   "
            This option specifies the test for the rmd algorithm"
    }
    cdl_component CYGPKG_OPENSSL_DES {
        display       "DES algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the DES Algorith."

        compile        crypto/des/set_key.c    \
                       crypto/des/ecb_enc.c    \
                       crypto/des/cbc_enc.c    \
                       crypto/des/ecb3_enc.c   \
                       crypto/des/cfb64enc.c   \
                       crypto/des/cfb64ede.c   \
                       crypto/des/cfb_enc.c    \
                       crypto/des/ofb64ede.c   \
                       crypto/des/enc_read.c   \
                       crypto/des/enc_writ.c   \
                       crypto/des/ofb64enc.c   \
                       crypto/des/ofb_enc.c    \
                       crypto/des/str2key.c    \
                       crypto/des/pcbc_enc.c   \
                       crypto/des/qud_cksm.c   \
                       crypto/des/rand_key.c   \
                       crypto/des/des_enc.c    \
                       crypto/des/fcrypt.c     \
                       crypto/des/fcrypt_b.c   \
                       crypto/des/xcbc_enc.c   \
                       crypto/des/rpc_enc.c    \
                       crypto/des/cbc_cksm.c   \
                       crypto/des/ede_cbcm_enc.c 

        cdl_component CYGPKG_OPENSSL_DES_READ_PWD {
            display       "DES read passwd from TTY"
            flavor        bool
            requires      CYGPKG_IO_SERIAL_TERMIOS
            requires      CYGPKG_IO_SERIAL_TERMIOS_TERMIOS0
            default_value 0
            description   "
                  Implement reading the passwd from the terminal.
                  This requires termios etc so is not compiled by
                  default. If you do use it make sure you have
                  termio0 correctly configured."

            compile   crypto/des/read2pwd.c   \
                      crypto/des/read_pwd.c   
        }               
    }                
    cdl_option CYGPKG_OPENSSL_DES_TESTS {
        display "OpenSSL DES tests"
        flavor  data
        no_define
        calculated { 
           " tests/destest.c"
        }
        description   "
            This option specifies the test for the DES algorithm"
    }
    cdl_option CYGPKG_OPENSSL_DES_READ_PWD_TESTS {
        display "OpenSSL DES read passwd tests"
        flavor data
        no_define
        calculated {
           " tests/despwdtest.c "
        }
        description   "
            This option specifies the test for the DES functions that
            read passwds from the user. The test it to ensure that 
            the passwd is not echoed."
    }
    cdl_component CYGPKG_OPENSSL_RC4 {
        display       "RC4 algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the RC4 Algorith."

        compile       crypto/rc4/rc4_skey.c   \
                      crypto/rc4/rc4_enc.c
    }                
    cdl_option CYGPKG_OPENSSL_RC4_TESTS {
        display "OpenSSL RC4 tests"
        flavor  data
        no_define
        calculated { 
           " tests/rc4test.c"
        }
        description   "
            This option specifies the test for the RC4 algorithm"
    }
    cdl_component CYGPKG_OPENSSL_RC2 {
        display       "RC2 algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the RC2 Algorith."

        compile        crypto/rc2/rc2_ecb.c    \
                       crypto/rc2/rc2_skey.c   \
                       crypto/rc2/rc2_cbc.c    \
                       crypto/rc2/rc2cfb64.c   \
                       crypto/rc2/rc2ofb64.c
    }                
    cdl_option CYGPKG_OPENSSL_RC2_TESTS {
        display "OpenSSL RC2 tests"
        flavor  data
        no_define
        calculated { 
           " tests/rc2test.c"
        }
        description   "
            This option specifies the test for the RC2 algorithm"
    }
    cdl_component CYGPKG_OPENSSL_BLOWFISH {
        display       "Blowfish algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the Blowfish Algorith."

        compile       crypto/bf/bf_skey.c     \
                      crypto/bf/bf_ecb.c      \
                      crypto/bf/bf_enc.c      \
                      crypto/bf/bf_cfb64.c    \
                      crypto/bf/bf_ofb64.c    

        cdl_option CYGPKG_OPENSSL_BLOWFISH_TESTS {
            display "OpenSSL Blowfist tests"
            flavor  data
            no_define
            calculated { 
               " tests/bftest.c"
            }
            description   "
                This option specifies the test for the Blowfish algorithm"
        }
    }
    cdl_component CYGPKG_OPENSSL_CAST {
        display       "Cast algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the Cast Algorith."

        compile       crypto/cast/c_skey.c    \
                      crypto/cast/c_ecb.c     \
                      crypto/cast/c_cfb64.c   \
                      crypto/cast/c_ofb64.c   \
                      crypto/cast/c_enc.c     

        cdl_option CYGPKG_OPENSSL_CAST_TESTS {
            display "OpenSSL Cast tests"
            flavor  data
            no_define
            calculated { 
               " tests/casttest.c"
            }
            description   "
                This option specifies the test for the CAST algorithm"
        }
    }
    cdl_component CYGPKG_OPENSSL_MDC2 {
        display       "MDC2 algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        requires      CYGPKG_OPENSSL_DES
        default_value 1
        description   "
             Implements the MDC2 Algorith."

        compile       crypto/mdc2/mdc2dgst.c  \
                      crypto/mdc2/mdc2_one.c 

        cdl_option CYGPKG_OPENSSL_MDC2_TESTS {
            display "OpenSSL MDC2 tests"
            flavor  data
            no_define
            calculated { 
               " tests/mdc2test.c"
            }
            description   "
                This option specifies the test for the MDC2 algorithm"
        }
    }
    cdl_component CYGPKG_OPENSSL_DSA {
        display       "DSA algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        requires      CYGPKG_OPENSSL_SHA1
        default_value 1
        description   "
             Implements the DSA Algorith."

        compile       crypto/dsa/dsa_gen.c    \
                      crypto/dsa/dsa_key.c    \
                      crypto/dsa/dsa_lib.c    \
                      crypto/dsa/dsa_asn1.c   \
                      crypto/dsa/dsa_vrf.c    \
                      crypto/dsa/dsa_sign.c   \
                      crypto/dsa/dsa_err.c    \
                      crypto/dsa/dsa_ossl.c   \

        cdl_option CYGPKG_OPENSSL_DSA_TESTS {
            display "OpenSSL DSA tests"
            flavor  data
            no_define
            calculated { 
               " tests/dsatest.c"
            }
            description   "
                This option specifies the test for the DSA algorithm"
        }
    }
    cdl_component CYGPKG_OPENSSL_DH {
        display       "DH algorithm"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the DH Algorith."

        compile        crypto/dh/dh_gen.c      \
                       crypto/dh/dh_key.c      \
                       crypto/dh/dh_lib.c      \
                       crypto/dh/dh_check.c    \
                       crypto/dh/dh_err.c     
    }
    cdl_option CYGPKG_OPENSSL_DH_TESTS {
        display "OpenSSL DH tests"
        flavor  data
        no_define
        calculated { 
           " tests/dhtest.c"
        }
        description   "
            This option specifies the test for the DH algorithm"
    }
    cdl_component CYGPKG_OPENSSL_BIO {
        display       "BIO API"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the BIO API"

        compile       crypto/bio/bio_lib.c    \
                      crypto/bio/bio_cb.c     \
                      crypto/bio/bio_err.c    \
                      crypto/bio/bss_mem.c    \
                      crypto/bio/bss_null.c   \
                      crypto/bio/bss_fd.c     \
                      crypto/bio/bss_file.c   \
                      crypto/bio/bss_sock.c   \
                      crypto/bio/bss_conn.c   \
                      crypto/bio/bf_null.c    \
                      crypto/bio/bf_buff.c    \
                      crypto/bio/b_print.c    \
                      crypto/bio/b_dump.c     \
                      crypto/bio/b_sock.c     \
                      crypto/bio/bss_acpt.c   \
                      crypto/bio/bf_nbio.c    \
                      crypto/bio/bss_log.c    \
                      crypto/bio/bss_bio.c    
    }
    cdl_component CYGPKG_OPENSSL_BUFFER {
        display       "Buffer API"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the buffer API"

        compile       crypto/buffer/buffer.c  \
                      crypto/buffer/buf_err.c 
    }

    cdl_component CYGPKG_OPENSSL_COMP {
        display       "COMP API"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the Compression API"

        compile       crypto/comp/comp_lib.c  \
                      crypto/comp/c_rle.c     \
                      crypto/comp/c_zlib.c    \
    }
    cdl_component CYGPKG_OPENSSL_ERR {
        display       "ERR API"
        flavor        bool
        requires      CYGPKG_OPENSSL
        default_value 1
        description   "
             Implements the Error message API."
    }
    cdl_component CYGPKG_OPENSSL_SSL {
        display       "SSL API"
        flavor        bool
        requires      CYGPKG_OPENSSL
        requires      CYGPKG_OPENSSL_MD5
        requires      CYGPKG_OPENSSL_RC4
        requires      CYGPKG_OPENSSL_RC2
        requires      CYGPKG_OPENSSL_IDEA
        requires      CYGPKG_OPENSSL_DES
        requires      CYGPKG_OPENSSL_SHA
        requires      CYGPKG_OPENSSL_COMP
        default_value 0
        description   "
             Implements the SSL API"

        compile       ssl/bio_ssl.c           \
                      ssl/s23_pkt.c           \
                      ssl/s2_lib.c            \
                      ssl/s3_both.c           \
                      ssl/s3_meth.c           \
                      ssl/ssl_asn1.c          \
                      ssl/ssl_err2.c          \
                      ssl/ssl_stat.c          \
                      ssl/t1_lib.c            \
                      ssl/s23_clnt.c          \
                      ssl/s23_srvr.c          \
                      ssl/s2_meth.c           \
                      ssl/s3_clnt.c           \
                      ssl/s3_pkt.c            \
                      ssl/ssl_cert.c          \
                      ssl/ssl_lib.c           \
                      ssl/ssl_txt.c           \
                      ssl/t1_meth.c           \
                      ssl/s23_lib.c           \
                      ssl/s2_clnt.c           \
                      ssl/s2_pkt.c            \
                      ssl/s3_enc.c            \
                      ssl/s3_srvr.c           \
                      ssl/ssl_ciph.c          \
                      ssl/ssl_rsa.c           \
                      ssl/t1_clnt.c           \
                      ssl/t1_srvr.c           \
                      ssl/s23_meth.c          \
                      ssl/s2_enc.c            \
                      ssl/s2_srvr.c           \
                      ssl/s3_lib.c            \
                      ssl/ssl_algs.c          \
                      ssl/ssl_err.c           \
                      ssl/ssl_sess.c          \
                      ssl/t1_enc.c
    }
    cdl_component CYGPKG_OPENSSL_OPTIONS {
        display "OpenSSL build options"
        flavor  none
	no_define

        cdl_option CYGPKG_OPENSSL_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS -I$(PREFIX)/include/openssl" }
            description   "
                This option modifies the set of compiler flags for
                building the OpenSSL package.
	        These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_OPENSSL_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "-Wstrict-prototypes" }
            description   "
                This option modifies the set of compiler flags for
                building the OpenSSL package. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_OPENSSL_TESTS {
            display    "List off all tests"
            flavor      data
            no_define
            calculated  {" tests/randtest.c tests/exptest.c \
                             tests/bntest.c tests/hmactest.c " . 
                             ( is_enabled(CYGPKG_OPENSSL_IDEA) ? 
                                  get_data(CYGPKG_OPENSSL_IDEA_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_RC5) ? 
                                  get_data(CYGPKG_OPENSSL_RC5_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_RSA) ? 
                                  get_data(CYGPKG_OPENSSL_RSA_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_MD2) ? 
                                  get_data(CYGPKG_OPENSSL_MD2_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_MD4) ? 
                                  get_data(CYGPKG_OPENSSL_MD4_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_MD5) ? 
                                  get_data(CYGPKG_OPENSSL_MD5_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_SHA) ? 
                                  get_data(CYGPKG_OPENSSL_SHA_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_SHA1) ? 
                                  get_data(CYGPKG_OPENSSL_SHA1_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_RMD160) ? 
                                  get_data(CYGPKG_OPENSSL_RMD160_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_DES_READ_PWD) ? 
                                  get_data(CYGPKG_OPENSSL_DES_READ_PWD_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_DES) ? 
                                  get_data(CYGPKG_OPENSSL_DES_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_RC4) ? 
                                  get_data(CYGPKG_OPENSSL_RC4_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_RC2) ? 
                                  get_data(CYGPKG_OPENSSL_RC2_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_BLOWFISH) ? 
                                  get_data(CYGPKG_OPENSSL_BLOWFISH_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_CAST) ? 
                                  get_data(CYGPKG_OPENSSL_CAST_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_MDC2) ? 
                                  get_data(CYGPKG_OPENSSL_MDC2_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_DSA) ? 
                                  get_data(CYGPKG_OPENSSL_DSA_TESTS) :
                                  " " ) .
                             ( is_enabled(CYGPKG_OPENSSL_DH) ? 
                                  get_data(CYGPKG_OPENSSL_DH_TESTS) :
                                  " " ) 
                        }
            description   "
                This option specifies the set of tests for the eCos 
                OpenSSL library. The tests that get compiled depends
                on which parts of the library are enabled"
        }
    }
}

# EOF openssl.cdl
